// Shift type.
parameter LSL = 0;
parameter LSR = 1;
parameter ASR = 2;
parameter ROR = 3;
parameter RORI = 4;
