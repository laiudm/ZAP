// Modes
parameter FIQ = 5'b10_001;
parameter IRQ = 5'b10_010;
parameter ABT = 5'b10_111;
parameter SVC = 5'b10_011;
parameter USR = 5'b10_000;
parameter SYS = 5'b11_111;
parameter UND = 5'b11_011;
