// Shift type.
parameter [1:0] LSL = 0;
parameter [1:0] LSR = 1;
parameter [1:0] ASR = 2;
parameter [1:0] ROR = 3;
parameter [2:0] RORI = 4;
