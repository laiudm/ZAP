`default_nettype none

module zap_alu_stage #(
        parameter PHY_REGS = 46,
        parameter SHIFT_OPS = 5,
        parameter ALU_OPS = 32
)
(
        // ============================================
        // Clock and reset.
        // ============================================
        input wire                         i_clk,
        input wire                         i_reset,

        // ============================================
        // From CPSR. ( I, F, T, Mode )
        // ============================================
        input wire  [31:0]                 i_cpsr_ff,
        input wire  [31:0]                 i_cpsr_nxt,

        // =============================================
        // Clear and Stall signals.
        // =============================================
        input wire                      i_clear_from_writeback, // | High Priority
        input wire                      i_data_stall,           // V Low Priority

        // =============================================
        // Inputs from shift.
        // =============================================
        input wire  [31:0]                 i_mem_srcdest_value_ff,
        input wire  [31:0]                 i_alu_source_value_ff, 
        input wire  [31:0]                 i_shifted_source_value_ff,
        input wire                         i_shift_carry_ff,
        input wire                         i_rrx_ff,
        input wire  [31:0]                 i_pc_plus_8_ff,
        input wire  [3:0]                  i_interrupt_vector_ff,       // { IRQ, FIQ, I-ABT, SWI }
        input wire  [$clog2(PHY_REGS)-1:0] i_mem_srcdest_index_ff,     
        input wire  [8:0]                  i_mem_magic_number_ff,       // {LOAD, STORE, ... }
        input wire  [3:0]                  i_condition_code_ff,
        input wire  [$clog2(PHY_REGS)-1:0] i_destination_index_ff,
        input wire  [$clog2(ALU_OPS):0]    i_alu_operation_ff,          // { OP, S }
        input wire  [$clog2(SHIFT_OPS)-1:0]o_shift_operation_ff,

        // ===========================================
        // Outputs
        // ===========================================
        output reg [31:0]                   o_alu_result_nxt,
        output reg [31:0]                   o_alu_result_ff,
        output reg [8:0]                    o_mem_magic_number_ff,      
        output reg                          o_dav_ff,
        output reg [31:0]                   o_pc_plus_8_ff,
        output reg [31:0]                   o_mem_address_ff,           // Memory addresss sent. 
        output reg                          o_clear_from_alu,
        output reg [31:0]                   o_pc_from_alu,
        output reg [$clog2(PHY_REGS)-1:0]   o_destination_index_ff,
        output reg [3:0]                    o_interrupt_vector_ff,
        output reg [$clog2(PHY_REGS)-1:0]   o_mem_srcdest_index_ff,
        output reg              [3:0]       o_interrupt_vector_ff
);

`include "cc.vh"
`include "regs.vh"
`include "opcodes.vh"

localparam N = 3;
localparam Z = 2;
localparam C = 1;
localparam V = 0;

reg [31:0] o_dav_nxt;
reg [3:0] flags_ff, flags_nxt;
reg [31:0] rm, rn;
reg [31:0] mem_address_nxt;

reg mem_load_ff,                     
mem_store_ff,
mem_pre_index_ff,                
mem_unsigned_byte_enable_ff,     
mem_signed_byte_enable_ff,       
mem_signed_halfword_enable_ff,
mem_unsigned_halfword_enable_ff,
mem_translate_ff,                
force_locked_access_ff;

always @*
begin
        rm = i_shifted_source_value_ff;
        rn = i_alu_source_value_ff;
end

always @*
{mem_load_ff,                     
mem_store_ff,
mem_pre_index_ff,                
mem_unsigned_byte_enable_ff,     
mem_signed_byte_enable_ff,       
mem_signed_halfword_enable_ff,
mem_unsigned_halfword_enable_ff,
mem_translate_ff,                
force_locked_access_ff} = i_mem_magic_number_ff;

// ===========================================
// Provides branch instructions.
// ===========================================
always @*
begin
        // This is interesting...

        if ( i_destination_index_ff == PHY_PC )
        begin
                o_clear_from_alu = 1'd1;
                o_pc_from_alu    = o_alu_result_nxt;
        end
        else
        begin
                o_clear_from_alu = 1'd0;
                o_pc_from_alu = 32'd0;
        end
end

// ==========================================
// This check can be done independently of
// others.
// ==========================================
always @*
        o_dav_nxt = is_cc_satisfied ( i_condition_code_ff, flags_ff );

always @ (posedge i_clk)
begin
        if ( i_reset )
        begin
                flags_ff <= 0;
                o_dav_ff <= 0;
        end
        else if ( i_clear_from_writeback )
        begin
                o_dav_ff <= 0;
                flags_ff <= i_cpsr_nxt;
        end
        else if ( i_data_stall )
        begin
                // Preserve values.
        end
        else
        begin
                o_alu_result_ff         <= o_alu_result_nxt;
                o_mem_magic_number_ff   <= i_mem_magic_number_ff;
                o_dav_ff                <= o_dav_nxt;                
                o_pc_plus_8_ff          <= i_pc_plus_8_ff;
                o_mem_address_ff        <= mem_address_nxt;
                o_destination_index_ff  <= i_destination_index_ff;
                flags_ff                <= o_dav_nxt ? flags_nxt : flags_ff;
                o_interrupt_vector_ff   <= i_interrupt_vector_ff;
                o_mem_srcdest_index_ff  <= i_mem_srcdest_index_ff;
                o_interrupt_vector_ff   <= i_interrupt_vector_ff;
        end
end

always @*
begin: blk1
        reg [31:0] rd;
        reg [$clog2(ALU_OPS):0]  opcode;

        opcode = i_alu_operation_ff;

       o_dav_nxt = is_cc_satisfied ( i_condition_code_ff, flags_ff );

        if (    opcode == AND || 
                opcode == EOR || 
                opcode == MOV || 
                opcode == MVN || 
                opcode == BIC || 
                opcode == ORR )
        begin
                {flags_nxt, rd} = process_logical_instructions ( rn, rm, flags_ff, opcode );
        end
        else if ( opcode == FMOV || opcode == MMOV )
        begin: blk2
                // =============================================================
                // Update ALU flags if needed. Also a fancy MOV instruction.
                // =============================================================
                // This is a special kind of MOV instruction that has mask bits
                // in ALU source.

                integer i;
                reg [31:0] exp_mask;

                flags_nxt = flags_ff;

                rd = {flags_ff, 4'd0, 8'd0, 8'd0, i_cpsr_ff[7:0]}; 
                exp_mask = {{8{rn[3]}},{8{rn[2]}},{8{rn[1]}},{8{rn[0]}}};

                for ( i=0;i<32;i=i+1 )
                begin
                        if ( exp_mask[i] )
                                rd[i] = rm[i];
                end                
        end
        begin
                {flags_nxt, rd} = process_arithmetic_instructions ( rn, rm, flags_ff, opcode );
        end

        // ==========================
        // Memory address.
        // ==========================
        if ( mem_pre_index_ff == 1 )
                mem_address_nxt = rn;  
        else
                mem_address_nxt = rd;

        o_alu_result_nxt = rd;
end

// ===============================================================
// Process logical instructions.
// ===============================================================
function [35:0] process_logical_instructions 
( input [31:0] rn, rm, input [3:0] flags, input [$clog2(ALU_OPS):0] op );
begin: blk2
        reg [31:0] rd;
        reg [3:0] flags_out;

        case(op >> 1)
        AND: rd = rn & rm;
        EOR: rd = rn ^ rm;
        BIC: rd = rn & ~(rm);
        MOV: rd = rm;
        MVN: rd = ~rm;
        ORR: rd = rn | rm;
        TST: rd = rn & rm;
        TEQ: rd = rn ^ rn;
        endcase           

        flags_out = flags;

        if ( rd == 0 && op[0] )
                flags_out[Z] = 1'd1;

        if ( rd[31] && op[0] )
                flags_out[N] = 1'd1;

        process_logical_instructions = {flags_out, rd};     
end
endfunction

// ===============================================================
// Process arithmetic instructions.
// ===============================================================
function [35:0] process_arithmetic_instructions 
( input [31:0] rn, rm, input [3:0] flags, input [$clog2(ALU_OPS):0] op );
begin: blk3
        reg [31:0] rd;
        reg n,z,c,v;
        reg [3:0] flags_out;

        case ( op >> 1 )
        ADD: {c,rd} = rn +  rm + 32'd0;
        ADC: {c,rd} = rn +  rm + flags[C];
        SUB: {c,rd} = rn + ~rm + 32'd1;
        RSB: {c,rd} = rn + ~rm + 32'd1;
        SBC: {c,rd} = rn + ~rm + !flags[C];
        RSC: {c,rd} = rm + ~rn + !flags[C];
        CMP: {c,rd} = rm + ~rn + 32'd0;
        CMN: {c,rd} = rm + ~rn + 32'd1;
        endcase

        flags_out = flags;

        if ( op[0] )
        begin
                if ( rd == 0 )                  flags_out[Z] = 1;
                if ( rd[31] )                   flags_out[N] = 1;
                if ( c )                        flags_out[C] = 1;

                // Overflow.
                if ( rn[31] == rm[31] && (rd[31] != rn[31]) )
                begin
                        flags_out[V] = 1;
                end 
        end

        process_arithmetic_instructions = {flags_out, rd};

end
endfunction

// ===============================================================
// Determines if the current instruction is worthy of execution.
// ===============================================================
function is_cc_satisfied 
( 
        input [3:0] cc,         // 31:28 of the instruction. 
        input [3:0] fl          // CPSR flags.
);
reg ok,n,z,c,v;
begin
        {n,z,c,v} = fl;

        case(cc)
        EQ:     ok =  z;
        NE:     ok = !z;
        CS:     ok = c;
        CC:     ok = !c;
        MI:     ok = n;
        PL:     ok = !n;
        VS:     ok = v;
        VC:     ok = !v;
        HI:     ok = c && !z;
        LS:     ok = !c || z;
        GE:     ok = n^v;
        LT:     ok = !(n^v);
        GT:     ok = (n^v) && !z;
        LE:     ok = (!(n^v)) || z;
        AL:     ok = 1;
        NV:     ok = 0;                    
        endcase   

        is_cc_satisfied = ok;
end
endfunction

endmodule
