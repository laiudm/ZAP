`ifndef __FIELDS_VH__
`define __FIELDS_VH__

`define BASE_EXTEND             33
`define BASE                    19:16
`define SRCDEST_EXTEND          32
`define SRCDEST                 15:12
`define DP_RD_EXTEND            33      // Destination source extend.
`define DP_RD                   15:12   // Destination source.
`define DP_RS_EXTEND            32      // Shift source extend.
`define DP_RS                   3:0     // Shift source. ARM refers to this as rm.
`define DP_RN                   19:16   // ALU source.
`define DP_RN_EXTEND            34      // ALU source extend.
`define OPCODE_EXTEND           35      // To differential lower and higher -> 1 means higher.

`endif
