//
// For transferring indices/immediates across stages.
//
parameter              INDEX_EN       =       1'd0;
parameter              IMMED_EN       =       1'd1;
