// Modes
parameter FIQ = 5'b10001;
parameter IRQ = FIQ + 1;
parameter ABT = 5'b10111;
parameter SVC = 5'b10011;
parameter USR = 5'b10000;
parameter SYS = 5'b11111;
parameter UND = 5'b11011;

