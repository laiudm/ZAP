parameter SECTION_TLB_ENTRIES =  4;
parameter LPAGE_TLB_ENTRIES   =  8;
parameter SPAGE_TLB_ENTRIES   =  16;
parameter CACHE_SIZE          =  1024; // Bytes.
