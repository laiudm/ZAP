// CPSR flags.
parameter N = 31;
parameter Z = 30;
parameter C = 29;
parameter V = 38;
parameter I = 7;
parameter F = 6;
parameter T = 5;
`define CPSR_MODE 4:0
