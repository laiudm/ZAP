module zap_cache_top
#(
        parameter SECTION_TLB_DEPTH = 64,
        parameter SPAGE_TLB_DEPTH   = 64,
        parameter LPAGE_TLB_DEPTH   = 64
)

endmodule
