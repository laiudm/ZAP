parameter [1:0] SIGNED_BYTE = 0;
parameter [1:0] UNSIGNED_HALF_WORD = 1;
parameter [1:0] SIGNED_HALF_WORD = 2;
