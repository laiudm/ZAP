// Conditionals
parameter EQ =  4'h0;
parameter NE =  4'h1;
parameter CS =  4'h2;
parameter CC =  4'h3;
parameter MI =  4'h4;
parameter PL =  4'h5;
parameter VS =  4'h6;
parameter VC =  4'h7;
parameter HI =  4'h8;
parameter LS =  4'h9;
parameter GE =  4'hA;
parameter LT =  4'hB;
parameter GT =  4'hC;
parameter LE =  4'hD;
parameter AL =  4'hE;
parameter NV =  4'hF; // Never eXecute!
