// CPSR flags.
parameter N = 31;
parameter Z = 30;
parameter C = 29;
parameter V = 38;
